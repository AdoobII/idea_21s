LIBRARY ieee;
USE ieee.numeric_std.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY idea IS
    PORT (
        X_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        X_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        X_3 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        X_4 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        KEY : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
        Y_1 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        Y_2 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        Y_3 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        Y_4 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END idea;

ARCHITECTURE Behavioral OF idea IS

    --  Component Declaration for ROUND, TRAFO
    --  ROUND
    COMPONENT round_module
        PORT (
            X_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_3 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_4 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_3 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_4 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_5 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_6 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_1 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_2 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_3 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_4 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
    END COMPONENT;
    --  TRAFO
    COMPONENT trafo
        PORT (
            X_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_3 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            X_4 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_3 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Z_4 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_1 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_2 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_3 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
            Y_4 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
    END COMPONENT;
    --KEYGEN
    COMPONENT keygen
        PORT (
            KEY : IN STD_LOGIC_VECTOR (127 DOWNTO 0);
            ROUND_KEY_1 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_2 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_3 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_4 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_5 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_6 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_7 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            ROUND_KEY_8 : OUT STD_LOGIC_VECTOR(95 DOWNTO 0);
            TRAFO_KEY_1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
        );
    END COMPONENT;

    --signals
    --round outputs
    SIGNAL ROUND_O_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    SIGNAL ROUND_O_8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
    --partial keys
    SIGNAL ROUND_KEY_1 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_2 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_3 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_4 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_5 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_6 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_7 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL ROUND_KEY_8 : STD_LOGIC_VECTOR(95 DOWNTO 0);
    SIGNAL TRAFO_KEY_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
BEGIN
    --INSTANTIATE KEYGEN TO GET THE 54 PARTIAL KEYS
    cKEYGEN_1 : keygen PORT MAP(
        KEY => KEY, ROUND_KEY_1 => ROUND_KEY_1, ROUND_KEY_2 => ROUND_KEY_2,
        ROUND_KEY_3 => ROUND_KEY_3, ROUND_KEY_4 => ROUND_KEY_4,
        ROUND_KEY_5 => ROUND_KEY_5, ROUND_KEY_6 => ROUND_KEY_6,
        ROUND_KEY_7 => ROUND_KEY_7, ROUND_KEY_8 => ROUND_KEY_8,
        TRAFO_KEY_1 => TRAFO_KEY_1);
    --Instantiate ROUND modules
    cROUND_1 : round_module PORT MAP(
        X_1, X_2, X_3, X_4,
        Z_1 => ROUND_KEY_1(95 DOWNTO 80), Z_2 => ROUND_KEY_1(79 DOWNTO 64),
        Z_3 => ROUND_KEY_1(63 DOWNTO 48), Z_4 => ROUND_KEY_1(47 DOWNTO 32),
        Z_5 => ROUND_KEY_1(31 DOWNTO 16), Z_6 => ROUND_KEY_1(15 DOWNTO 0),
        Y_1 => ROUND_O_1(63 DOWNTO 48), Y_2 => ROUND_O_1(47 DOWNTO 32),
        Y_3 => ROUND_O_1(31 DOWNTO 16), Y_4 => ROUND_O_1(15 DOWNTO 0));

    cROUND_2 : round_module PORT MAP(
        X_1 => ROUND_O_1(63 DOWNTO 48), X_2 => ROUND_O_1(47 DOWNTO 32),
        X_3 => ROUND_O_1(31 DOWNTO 16), X_4 => ROUND_O_1(15 DOWNTO 0),
        Z_1 => ROUND_KEY_2(95 DOWNTO 80), Z_2 => ROUND_KEY_2(79 DOWNTO 64),
        Z_3 => ROUND_KEY_2(63 DOWNTO 48), Z_4 => ROUND_KEY_2(47 DOWNTO 32),
        Z_5 => ROUND_KEY_2(31 DOWNTO 16), Z_6 => ROUND_KEY_2(15 DOWNTO 0),
        Y_1 => ROUND_O_2(63 DOWNTO 48), Y_2 => ROUND_O_2(47 DOWNTO 32),
        Y_3 => ROUND_O_2(31 DOWNTO 16), Y_4 => ROUND_O_2(15 DOWNTO 0));

    cROUND_3 : round_module PORT MAP(
        X_1 => ROUND_O_2(63 DOWNTO 48), X_2 => ROUND_O_2(47 DOWNTO 32),
        X_3 => ROUND_O_2(31 DOWNTO 16), X_4 => ROUND_O_2(15 DOWNTO 0),
        Z_1 => ROUND_KEY_3(95 DOWNTO 80), Z_2 => ROUND_KEY_3(79 DOWNTO 64),
        Z_3 => ROUND_KEY_3(63 DOWNTO 48), Z_4 => ROUND_KEY_3(47 DOWNTO 32),
        Z_5 => ROUND_KEY_3(31 DOWNTO 16), Z_6 => ROUND_KEY_3(15 DOWNTO 0),
        Y_1 => ROUND_O_3(63 DOWNTO 48), Y_2 => ROUND_O_3(47 DOWNTO 32),
        Y_3 => ROUND_O_3(31 DOWNTO 16), Y_4 => ROUND_O_3(15 DOWNTO 0));

    cROUND_4 : round_module PORT MAP(
        X_1 => ROUND_O_3(63 DOWNTO 48), X_2 => ROUND_O_3(47 DOWNTO 32),
        X_3 => ROUND_O_3(31 DOWNTO 16), X_4 => ROUND_O_3(15 DOWNTO 0),
        Z_1 => ROUND_KEY_4(95 DOWNTO 80), Z_2 => ROUND_KEY_4(79 DOWNTO 64),
        Z_3 => ROUND_KEY_4(63 DOWNTO 48), Z_4 => ROUND_KEY_4(47 DOWNTO 32),
        Z_5 => ROUND_KEY_4(31 DOWNTO 16), Z_6 => ROUND_KEY_4(15 DOWNTO 0),
        Y_1 => ROUND_O_4(63 DOWNTO 48), Y_2 => ROUND_O_4(47 DOWNTO 32),
        Y_3 => ROUND_O_4(31 DOWNTO 16), Y_4 => ROUND_O_4(15 DOWNTO 0));

    cROUND_5 : round_module PORT MAP(
        X_1 => ROUND_O_4(63 DOWNTO 48), X_2 => ROUND_O_4(47 DOWNTO 32),
        X_3 => ROUND_O_4(31 DOWNTO 16), X_4 => ROUND_O_4(15 DOWNTO 0),
        Z_1 => ROUND_KEY_5(95 DOWNTO 80), Z_2 => ROUND_KEY_5(79 DOWNTO 64),
        Z_3 => ROUND_KEY_5(63 DOWNTO 48), Z_4 => ROUND_KEY_5(47 DOWNTO 32),
        Z_5 => ROUND_KEY_5(31 DOWNTO 16), Z_6 => ROUND_KEY_5(15 DOWNTO 0),
        Y_1 => ROUND_O_5(63 DOWNTO 48), Y_2 => ROUND_O_5(47 DOWNTO 32),
        Y_3 => ROUND_O_5(31 DOWNTO 16), Y_4 => ROUND_O_5(15 DOWNTO 0));

    cROUND_6 : round_module PORT MAP(
        X_1 => ROUND_O_5(63 DOWNTO 48), X_2 => ROUND_O_5(47 DOWNTO 32),
        X_3 => ROUND_O_5(31 DOWNTO 16), X_4 => ROUND_O_5(15 DOWNTO 0),
        Z_1 => ROUND_KEY_6(95 DOWNTO 80), Z_2 => ROUND_KEY_6(79 DOWNTO 64),
        Z_3 => ROUND_KEY_6(63 DOWNTO 48), Z_4 => ROUND_KEY_6(47 DOWNTO 32),
        Z_5 => ROUND_KEY_6(31 DOWNTO 16), Z_6 => ROUND_KEY_6(15 DOWNTO 0),
        Y_1 => ROUND_O_6(63 DOWNTO 48), Y_2 => ROUND_O_6(47 DOWNTO 32),
        Y_3 => ROUND_O_6(31 DOWNTO 16), Y_4 => ROUND_O_6(15 DOWNTO 0));

    cROUND_7 : round_module PORT MAP(
        X_1 => ROUND_O_6(63 DOWNTO 48), X_2 => ROUND_O_6(47 DOWNTO 32),
        X_3 => ROUND_O_6(31 DOWNTO 16), X_4 => ROUND_O_6(15 DOWNTO 0),
        Z_1 => ROUND_KEY_7(95 DOWNTO 80), Z_2 => ROUND_KEY_7(79 DOWNTO 64),
        Z_3 => ROUND_KEY_7(63 DOWNTO 48), Z_4 => ROUND_KEY_7(47 DOWNTO 32),
        Z_5 => ROUND_KEY_7(31 DOWNTO 16), Z_6 => ROUND_KEY_7(15 DOWNTO 0),
        Y_1 => ROUND_O_7(63 DOWNTO 48), Y_2 => ROUND_O_7(47 DOWNTO 32),
        Y_3 => ROUND_O_7(31 DOWNTO 16), Y_4 => ROUND_O_7(15 DOWNTO 0));

    cROUND_8 : round_module PORT MAP(
        X_1 => ROUND_O_7(63 DOWNTO 48), X_2 => ROUND_O_7(47 DOWNTO 32),
        X_3 => ROUND_O_7(31 DOWNTO 16), X_4 => ROUND_O_7(15 DOWNTO 0),
        Z_1 => ROUND_KEY_8(95 DOWNTO 80), Z_2 => ROUND_KEY_8(79 DOWNTO 64),
        Z_3 => ROUND_KEY_8(63 DOWNTO 48), Z_4 => ROUND_KEY_8(47 DOWNTO 32),
        Z_5 => ROUND_KEY_8(31 DOWNTO 16), Z_6 => ROUND_KEY_8(15 DOWNTO 0),
        Y_1 => ROUND_O_8(63 DOWNTO 48), Y_2 => ROUND_O_8(47 DOWNTO 32),
        Y_3 => ROUND_O_8(31 DOWNTO 16), Y_4 => ROUND_O_8(15 DOWNTO 0));

    --Instantiate TRAFO
    cTRAFO_1 : trafo PORT MAP(
        X_1 => ROUND_O_8(63 DOWNTO 48), X_2 => ROUND_O_8(47 DOWNTO 32),
        X_3 => ROUND_O_8(31 DOWNTO 16), X_4 => ROUND_O_8(15 DOWNTO 0),
        Z_1 => TRAFO_KEY_1(63 DOWNTO 48), Z_2 => TRAFO_KEY_1(47 DOWNTO 32),
        Z_3 => TRAFO_KEY_1(31 DOWNTO 16), Z_4 => TRAFO_KEY_1(15 DOWNTO 0),
        Y_1 => Y_1, Y_2 => Y_2, Y_3 => Y_3, Y_4 => Y_4);
END Behavioral;