LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY xorop IS
	PORT (
		I_1 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		I_2 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		O_1 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END xorop;

ARCHITECTURE Behavioral OF xorop IS

BEGIN

	XOROP_proc : PROCESS (I_1, I_2)
	BEGIN
		O_1 <= (I_1 XOR I_2);
	END PROCESS XOROP_proc;

END Behavioral;